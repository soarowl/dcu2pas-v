module main

interface IDecoder {
	decode() !
	int_str() string
	imp_str() string
}
