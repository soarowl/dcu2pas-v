module main

interface IDecoder {
	int_str() string
	imp_str() string
}
